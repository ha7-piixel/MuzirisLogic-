//Verilog module for Muziris Logic
module Muziris_Gate(input wire a, input wire b, output wire y);
	assign y = a & b;
endmodule
